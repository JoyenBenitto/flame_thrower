package crossbar;


endpackage crossbar