/*
Idea is to use bluecheck to create synthesizable testbench
*/